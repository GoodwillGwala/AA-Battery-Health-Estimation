* LMX24_LM2902 - Rev. A
* Created by Paul Goedeke; November 16, 2018
* Created with Green-Williams-Lis Op Amp Macro-model Architecture
* Copyright 2018 by Texas Instruments Corporation
******************************************************
* MACRO-MODEL SIMULATED PARAMETERS:
******************************************************
* OPEN-LOOP GAIN AND PHASE VS. FREQUENCY  WITH RL, CL EFFECTS (Aol)
* UNITY GAIN BANDWIDTH (GBW)
* INPUT COMMON-MODE REJECTION RATIO VS. FREQUENCY (CMRR)
* POWER SUPPLY REJECTION RATIO VS. FREQUENCY (PSRR)
* DIFFERENTIAL INPUT IMPEDANCE (Zid)
* COMMON-MODE INPUT IMPEDANCE (Zic)
* OPEN-LOOP OUTPUT IMPEDANCE VS. FREQUENCY (Zo)
* OUTPUT CURRENT THROUGH THE SUPPLY (Iout)
* INPUT VOLTAGE NOISE DENSITY VS. FREQUENCY (en)
* INPUT CURRENT NOISE DENSITY VS. FREQUENCY (in)
* OUTPUT VOLTAGE SWING vs. OUTPUT CURRENT (Vo)
* SHORT-CIRCUIT OUTPUT CURRENT (Isc)
* QUIESCENT CURRENT (Iq)
* SETTLING TIME VS. CAPACITIVE LOAD (ts)
* SLEW RATE (SR)
* SMALL SIGNAL OVERSHOOT VS. CAPACITIVE LOAD
* LARGE SIGNAL RESPONSE
* OVERLOAD RECOVERY TIME (tor)
* INPUT BIAS CURRENT (Ib)
* INPUT OFFSET CURRENT (Ios)
* INPUT OFFSET VOLTAGE (Vos)
* INPUT COMMON-MODE VOLTAGE RANGE (Vcm)
* INPUT OFFSET VOLTAGE VS. INPUT COMMON-MODE VOLTAGE (Vos vs. Vcm)
* INPUT/OUTPUT ESD CELLS (ESDin, ESDout)
******************************************************
.subckt LMX24_LM2902 IN+ IN- VCC VEE OUT
******************************************************
* MODEL DEFINITIONS:
.model BB_SW VSWITCH(Ron=50 Roff=1e12 Von=700e-3 Voff=0)
.model ESD_SW VSWITCH(Ron=50 Roff=1e12 Von=250e-3 Voff=0)
.model OL_SW VSWITCH(Ron=1e-3 Roff=1e9 Von=900e-3 Voff=800e-3)
.model OR_SW VSWITCH(Ron=10e-3 Roff=1e9 Von=1e-3 Voff=0)
.model R_NOISELESS RES(T_ABS=-273.15)
******************************************************


I_OS        ESDn MID -18N
I_B         37 MID -20N
V_GRp       57 MID 180
V_GRn       58 MID -180
V_ISCp      51 MID 40
V_ISCn      52 MID -40
V_ORn       45 VCLP -1.2
V11         56 44 0
V_ORp       43 VCLP 1.2
V12         55 42 0
V4          33 OUT 0
VCM_MIN     79 VEE_B 0
VCM_MAX     80 VCC_B -1.5
I_Q         VCC VEE 175U
V_OS        86 37 1.8M
R61         MID 22 R_NOISELESS 8.001K 
C16         22 23 19.89P 
R58         23 22 R_NOISELESS 100MEG 
GVCCS2      23 MID VEE_B MID  -992.9M
R57         MID 23 R_NOISELESS 1 
XU3         VCC_B VEE_B 24 25 26 27 MID PHASEREV_0
XU1         VIMON MID CRS CRS_DIST_0
C21         28 29 313.8N  
C22         30 31 636.6F  
R70         31 MID R_NOISELESS 2.5 
R67         31 30 R_NOISELESS 10K 
R66         30 MID R_NOISELESS 1 
XU2         31 MID MID 32 VCCS_LIM_ZO_0
GVCCS4      30 MID 29 MID  -4.3
R65         29 MID R_NOISELESS 3.03K 
R64         29 28 R_NOISELESS 10K 
R63         28 MID R_NOISELESS 1 
GVCCS3      28 MID CL_CLAMP 33  -90
R62         32 MID R_NOISELESS 1 
C29         34 MID 47F 
R78         MID 34 R_NOISELESS 1MEG 
GVCCS9      34 MID 35 MID  -1U
XU5         36 MID MID CLAMP CRS MID VCCS_LIM_2_EN_0
C28         38 MID 1P 
R77         39 38 R_NOISELESS 100 
C27         40 MID 1P 
R76         41 40 R_NOISELESS 100 
R75         MID 42 R_NOISELESS 1 
GVCCS8      42 MID 43 MID  -1
R74         44 MID R_NOISELESS 1 
GVCCS7      44 MID 45 MID  -1
Xi_nn       ESDn MID FEMT_0
Xi_np       MID 37 FEMT_0
Xe_n        ESDp 37 VNSE_0
C25         35 MID 47F 
R69         MID 35 R_NOISELESS 1MEG 
GVCCS6      35 MID VSENSE MID  -1U
C20         CLAMP MID 9N 
R68         MID CLAMP R_NOISELESS 1MEG 
R44         MID 36 R_NOISELESS 1MEG 
XVCCS_LIM_1 46 27 MID 36 VCCS_LIM_1_0
Rdummy      MID 33 R_NOISELESS 25K 
Rx          33 32 R_NOISELESS 250K 
R56         MID 47 R_NOISELESS 1K 
C15         47 48 1.592P 
R55         48 47 R_NOISELESS 100MEG 
GVCCS1      48 MID VCC_B MID  -100M
R54         MID 48 R_NOISELESS 1 
R49         MID 49 R_NOISELESS 4.616K 
C14         49 50 26.53P 
R48         50 49 R_NOISELESS 100MEG 
G_adjust    50 MID ESDp MID  -685.2M
Rsrc        MID 50 R_NOISELESS 1 
XIQPos      VIMON MID MID VCC VCCS_LIMIT_IQ_0
XIQNeg      MID VIMON VEE MID VCCS_LIMIT_IQ_0
C_DIFF      ESDp ESDn 1P 
XCL_AMP     51 52 VIMON MID 53 54 CLAMP_AMP_LO_0
SOR_SWp     CLAMP 55 CLAMP 55  S_VSWITCH_1
SOR_SWn     56 CLAMP 56 CLAMP  S_VSWITCH_2
XGR_AMP     57 58 59 MID 60 61 CLAMP_AMP_HI_0
R39         57 MID R_NOISELESS 1T 
R37         58 MID R_NOISELESS 1T 
R42         VSENSE 59 R_NOISELESS 1M 
C19         59 MID 1F 
R38         60 MID R_NOISELESS 1 
R36         MID 61 R_NOISELESS 1 
R40         60 62 R_NOISELESS 1M 
R41         61 63 R_NOISELESS 1M 
C17         62 MID 1F 
C18         MID 63 1F 
XGR_SRC     62 63 CLAMP MID VCCS_LIM_GR_0
R21         53 MID R_NOISELESS 1 
R20         MID 54 R_NOISELESS 1 
R29         53 64 R_NOISELESS 1M 
R30         54 65 R_NOISELESS 1M 
C9          64 MID 1F 
C8          MID 65 1F 
XCL_SRC     64 65 CL_CLAMP MID VCCS_LIM_4_0
R22         51 MID R_NOISELESS 1T 
R19         MID 52 R_NOISELESS 1T 
XCLAWp      VIMON MID 66 VCC_B VCCS_LIM_CLAW+_0
XCLAWn      MID VIMON VEE_B 67 VCCS_LIM_CLAW-_0
R12         66 VCC_B R_NOISELESS 1K 
R16         66 68 R_NOISELESS 1M 
R13         VEE_B 67 R_NOISELESS 1K 
R17         69 67 R_NOISELESS 1M 
C6          69 MID 1F 
C5          MID 68 1F 
G2          VCC_CLP MID 68 MID  -1M
R15         VCC_CLP MID R_NOISELESS 1K 
G3          VEE_CLP MID 69 MID  -1M
R14         MID VEE_CLP R_NOISELESS 1K 
XCLAW_AMP   VCC_CLP VEE_CLP VOUT_S MID 70 71 CLAMP_AMP_LO_0
R26         VCC_CLP MID R_NOISELESS 1T 
R23         VEE_CLP MID R_NOISELESS 1T 
R25         70 MID R_NOISELESS 1 
R24         MID 71 R_NOISELESS 1 
R27         70 72 R_NOISELESS 1M 
R28         71 73 R_NOISELESS 1M 
C11         72 MID 1F 
C10         MID 73 1F 
XCLAW_SRC   72 73 CLAW_CLAMP MID VCCS_LIM_3_0
H2          41 MID V11 -1
H3          39 MID V12 1
C12         SW_OL MID 100P 
R32         74 SW_OL R_NOISELESS 100 
R31         74 MID R_NOISELESS 1 
XOL_SENSE   MID 74 40 38 OL_SENSE_0
S1          28 29 SW_OL MID  S_VSWITCH_3
H1          75 MID V4 1K
S7          VEE OUT VEE OUT  S_VSWITCH_4
S6          OUT VCC OUT VCC  S_VSWITCH_5
R11         MID 76 R_NOISELESS 1T 
R18         76 VOUT_S R_NOISELESS 100 
C7          VOUT_S MID 10P 
E5          76 MID OUT MID  1
C13         VIMON MID 10P 
R33         75 VIMON R_NOISELESS 100 
R10         MID 75 R_NOISELESS 1T 
R47         77 VCLP R_NOISELESS 100 
C24         VCLP MID 100P 
E4          77 MID CL_CLAMP MID  1
R46         MID CL_CLAMP R_NOISELESS 1K 
G9          CL_CLAMP MID CLAW_CLAMP MID  -1M
R45         MID CLAW_CLAMP R_NOISELESS 1K 
G8          CLAW_CLAMP MID 34 MID  -1M
R43         MID VSENSE R_NOISELESS 1K 
G15         VSENSE MID CLAMP MID  -1M
C4          46 MID 1F 
R9          46 78 R_NOISELESS 1M 
R7          MID 79 R_NOISELESS 1T 
R6          80 MID R_NOISELESS 1T 
R8          MID 78 R_NOISELESS 1 
XVCM_CLAMP  26 MID 78 MID 80 79 VCCS_EXT_LIM_0
E1          MID 0 81 0  1
R89         VEE_B 0 R_NOISELESS 1 
R5          82 VEE_B R_NOISELESS 1M 
C3          82 0 1F 
R60         81 82 R_NOISELESS 1MEG 
C1          81 0 1 
R3          81 0 R_NOISELESS 1T 
R59         83 81 R_NOISELESS 1MEG 
C2          83 0 1F 
R4          VCC_B 83 R_NOISELESS 1M 
R88         VCC_B 0 R_NOISELESS 1 
G17         VEE_B 0 VEE 0  -1
G16         VCC_B 0 VCC 0  -1
R_PSR       84 24 R_NOISELESS 1K 
G_PSR       24 84 47 22  -1M
R2          25 ESDn R_NOISELESS 1M 
R1          84 85 R_NOISELESS 1M 
R_CMR       86 85 R_NOISELESS 1K 
G_CMR       85 86 49 MID  -1M
C_CMn       ESDn MID 2P 
C_CMp       MID ESDp 2P 
R53         ESDn MID R_NOISELESS 1T 
R52         MID ESDp R_NOISELESS 1T 
R35         IN- ESDn R_NOISELESS 10M 
R34         IN+ ESDp R_NOISELESS 10M 

.MODEL S_VSWITCH_1 VSWITCH (RON=10M ROFF=1T VON=10M VOFF=0)
.MODEL S_VSWITCH_2 VSWITCH (RON=10M ROFF=1T VON=10M VOFF=0)
.MODEL S_VSWITCH_3 VSWITCH (RON=1M ROFF=1T VON=500M VOFF=100M)
.MODEL S_VSWITCH_4 VSWITCH (RON=50 ROFF=1T VON=500M VOFF=450M)
.MODEL S_VSWITCH_5 VSWITCH (RON=50 ROFF=1T VON=500M VOFF=450M)

*.ENDS LMX24_LM2902
*
.SUBCKT PHASEREV_0  VCC VEE VIN+ VIN- VOUT+ VOUT- MID
E1 VOUT+ MID VALUE={IF(V(VIN+,MID)<V(VEE,MID)-0.3,V(VCC,MID),V(VIN+,MID))}
E2 VOUT- MID VALUE={IF(V(VIN-,MID)<V(VEE,MID)-0.3,V(VCC,MID),V(VIN-,MID))}
.ENDS
*


.SUBCKT CRS_DIST_0  VIMON MID OUT
V1 VREF MID -40M
ESHF VSHF MID VIMON VREF 1
GZC MID ZC VALUE = {SGN(V(VSHF,MID))}
R1 ZC MID 1
C1 ZC MID 2U
GCR MID OUT VALUE = {IF((ABS(V(ZC,MID))<=0.9),0,1)}
R2 OUT MID 1
.ENDS
*


.SUBCKT VCCS_LIM_ZO_0  VC+ VC- IOUT+ IOUT-
.PARAM GAIN = 4E3
.PARAM IPOS = 1E6
.PARAM INEG = -1E6
G1 IOUT+ IOUT- VALUE={LIMIT(GAIN*V(VC+,VC-),INEG,IPOS)}
.ENDS
*


.SUBCKT VCCS_LIM_2_EN_0  VC+ VC- IOUT+ IOUT- EN MID
.PARAM GAIN = 8.4E-4
.PARAM IPOS = 0.0048
.PARAM INEG = -0.0048
G1 IOUT+ IOUT- VALUE={LIMIT(GAIN*V(EN,MID)*V(VC+,VC-),INEG,IPOS)}
.ENDS
*


.SUBCKT FEMT_0  1 2
.PARAM FLWF=1E-3
.PARAM NLFF=500
.PARAM NVRF=500
.PARAM GLFF={PWR(FLWF,0.25)*NLFF/1164}
.PARAM RNVF={1.184*PWR(NVRF,2)}
.MODEL DVNF D KF={PWR(FLWF,0.5)/1E11} IS=1.0E-16
I1 0 7 10E-3
I2 0 8 10E-3
D1 7 0 DVNF
D2 8 0 DVNF
E1 3 6 7 8 {GLFF}
R1 3 0 1E9
R2 3 0 1E9
R3 3 6 1E9
E2 6 4 5 0 10
R4 5 0 {RNVF}
R5 5 0 {RNVF}
R6 3 4 1E9
R7 4 0 1E9
G1 1 2 3 4 1E-6
.ENDS
*


.SUBCKT VNSE_0  1 2
.PARAM FLW=10
.PARAM NLF=80
.PARAM NVR=35
.PARAM GLF={PWR(FLW,0.25)*NLF/1164}
.PARAM RNV={1.184*PWR(NVR,2)}
.MODEL DVN D KF={PWR(FLW,0.5)/1E11} IS=1.0E-16
I1 0 7 10E-3
I2 0 8 10E-3
D1 7 0 DVN
D2 8 0 DVN
E1 3 6 7 8 {GLF}
R1 3 0 1E9
R2 3 0 1E9
R3 3 6 1E9
E2 6 4 5 0 10
R4 5 0 {RNV}
R5 5 0 {RNV}
R6 3 4 1E9
R7 4 0 1E9
E3 1 2 3 4 1
.ENDS
*


.SUBCKT VCCS_LIM_1_0  VC+ VC- IOUT+ IOUT-
.PARAM GAIN = 1E-4
.PARAM IPOS = .5
.PARAM INEG = -.5
G1 IOUT+ IOUT- VALUE={LIMIT(GAIN*V(VC+,VC-),INEG,IPOS)}
.ENDS
*


.SUBCKT VCCS_LIMIT_IQ_0  VC+ VC- IOUT+ IOUT-
.PARAM GAIN = 1E-3
G1 IOUT- IOUT+ VALUE={IF( (V(VC+,VC-)<=0),0,GAIN*V(VC+,VC-) )}
.ENDS
*


.SUBCKT CLAMP_AMP_LO_0  VC+ VC- VIN COM VO+ VO-
.PARAM G=1
GVO+ COM VO+ VALUE = {IF(V(VIN,COM)>V(VC+,COM),((V(VIN,COM)-V(VC+,COM))*G),0)}
GVO- COM VO- VALUE = {IF(V(VIN,COM)<V(VC-,COM),((V(VC-,COM)-V(VIN,COM))*G),0)}
.ENDS
*


.SUBCKT CLAMP_AMP_HI_0  VC+ VC- VIN COM VO+ VO-
.PARAM G=10
GVO+ COM VO+ VALUE = {IF(V(VIN,COM)>V(VC+,COM),((V(VIN,COM)-V(VC+,COM))*G),0)}
GVO- COM VO- VALUE = {IF(V(VIN,COM)<V(VC-,COM),((V(VC-,COM)-V(VIN,COM))*G),0)}
.ENDS
*


.SUBCKT VCCS_LIM_GR_0  VC+ VC- IOUT+ IOUT-
.PARAM GAIN = 1
.PARAM IPOS = 0.013
.PARAM INEG = -0.013
G1 IOUT+ IOUT- VALUE={LIMIT(GAIN*V(VC+,VC-),INEG,IPOS)}
.ENDS
*


.SUBCKT VCCS_LIM_4_0  VC+ VC- IOUT+ IOUT-
.PARAM GAIN = 1
.PARAM IPOS = 1.04
.PARAM INEG = -1.04
G1 IOUT+ IOUT- VALUE={LIMIT(GAIN*V(VC+,VC-),INEG,IPOS)}
.ENDS
*


.SUBCKT VCCS_LIM_CLAW+_0  VC+ VC- IOUT+ IOUT-
G1 IOUT+ IOUT- TABLE {ABS(V(VC+,VC-))} =
+(0, 1.17E-03)
+(0.0046251, 1.17E-3)
+(0.15716, 1.21E-3)
+(1.3309, 1.28E-3)
+(35.075, 2.12E-3)
+(35.680, 2.55E-3)
+(36.033, 2.84E-3)
+(37.416, 7.97E-3)
.ENDS
*


.SUBCKT VCCS_LIM_CLAW-_0  VC+ VC- IOUT+ IOUT-
G1 IOUT+ IOUT- TABLE {ABS(V(VC+,VC-))} =
+(0.010, 2.50E-5)
+(0.070, 2.50E-5)
+(0.090, 5.80E-4)
+(0.100, 6.06E-4)
+(0.760, 7.14E-4) 
+(1.440, 7.62E-4)
+(8.000, 1.10E-3)
+(13.60, 1.55E-3)
+(15.45, 1.75E-3)
+(17.26, 2.15E-3)
+(18.87, 2.94E-3)
+(21.58, 4.50E-3)
+(25.53, 1.02E-2)
.ENDS
*



.SUBCKT VCCS_LIM_3_0  VC+ VC- IOUT+ IOUT-
.PARAM GAIN = 1
.PARAM IPOS = 0.435
.PARAM INEG = -0.435
G1 IOUT+ IOUT- VALUE={LIMIT(GAIN*V(VC+,VC-),INEG,IPOS)}
.ENDS
*


.SUBCKT OL_SENSE_0  COM SW+ OLN  OLP
GSW+ COM SW+ VALUE = {IF((V(OLN,COM)>10E-3 | V(OLP,COM)>10E-3),1,0)}
.ENDS
*


.SUBCKT VCCS_EXT_LIM_0  VIN+ VIN- IOUT- IOUT+ VP+ VP-
.PARAM GAIN = 1
G1 IOUT+ IOUT- VALUE={LIMIT(GAIN*V(VIN+,VIN-),V(VP-,VIN-), V(VP+,VIN-))}
.ENDS
*


.ENDS LMX24_LM2902


